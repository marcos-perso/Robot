/share/Projects/uSoC/design/synthesis/uSoCGenerators/DualRAM_8x32.vhd