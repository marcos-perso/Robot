/share/Projects/uSoC/design/synthesis/uSoCGenerators/ClockSynthesizer.vhd