/share/Projects/uSoC/design/synthesis/uSoCGenerators/RAM1024x32.vhd